library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use STD.textio.all; 
use IEEE.std_logic_textio.all;

entity Tea is
    port (
        clk             : in std_logic;
        enable          : in std_logic;
        vi              : in std_logic_vector (63 downto 0);
		  key             : in std_logic_vector(127 downto 0);
		  mode            : in std_logic;
		  reset				: in std_logic;
		  vo       	      : out std_logic_vector (63 downto 0)
	 );
end entity Tea;

architecture behave of Tea is

	component TeaCore is
		 port (
		     clk				: in std_logic;
			  mode			: in std_logic; 								-- 0 code 1 decode
			  key          : in std_logic_vector(127 downto 0);	-- key
		     vi      	   : in std_logic_vector (63 downto 0); 	-- input data
			  enable			: in std_logic;
		     vo      	   : out std_logic_vector (63 downto 0);	-- data output
		     ready 			: out std_logic 
		 );
	end component;
	
	component Arc4_Cypher is
		 port (
			  clk				   : in std_logic;
			  key             : in std_logic_vector(127 downto 0);	-- key
			  i_stream			: in std_logic_vector(31 downto 0);
			  o_stream			: out std_logic_vector(31 downto 0);
			  reset				: in std_logic;
			  out_ok				: out std_logic
		 );
	end component;
	
	component Arc4_Ksa is
	 port (
		  clk					: in std_logic;
		  key             : in std_logic_vector(127 downto 0);
		  reset				: in std_logic;
		  status				: out std_logic_vector(2047 downto 0);
		  ready				: out std_logic
	 );
	end component;
	
	signal round				: unsigned(5 downto 0) := "000000";
	
	signal s_vi					: std_logic_vector(63 downto 0);
	signal s_mode				: std_logic;
	signal s_key				: std_logic_vector(127 downto 0);
	signal s_vo					: std_logic_vector(63 downto 0);
	
	signal s_enable			: std_logic;
	signal s_ready_tea		: std_logic;
	
	signal s_arc4_key			:std_logic_vector(127 downto 0);
	signal s_arc4_i 			:std_logic_vector(31 downto 0);
	signal s_arc4_o 			:std_logic_vector(31 downto 0);
	
	signal s_key2      	  : std_logic_vector (127 downto 0);
	signal s_status		  : std_logic_vector(2047 downto 0);
	signal s_ready_arc	  : std_logic;
	signal s_out_ok		  : std_logic;
	
begin
	
	core1: TeaCore port map (
		clk => clk,
		mode => mode,
		key => key,
		vi => s_vi,		
		vo => s_vo,
		enable => s_enable,
		ready => s_ready_tea
	);
	
	arc4_1: Arc4_Cypher port map (
		clk => clk,
		key 		=> s_arc4_key,
	   i_stream	=> s_arc4_i,
		o_stream	=> s_arc4_o,
		reset => reset,
		out_ok => s_out_ok
	);
	
	Arc_i2 : Arc4_Ksa
        port map(
		      clk => clk,
				key 	 => s_key2,
				status => s_status,
				reset	=> reset,
				ready => s_ready_arc
    );
	
	process (clk, vi, s_vo) 
		variable mline : line;
	begin
	
		if(rising_edge(clk)) then
			
			if (enable = '1') then
			
				s_enable <= '1';
				
				if (round = "000000") then
						s_vi <= vi;
				elsif (round = "100000") then
						s_enable <= '0';
						vo <= s_vo;
				else 		
						s_vi <= s_vo;
				end if;
				
				round <= round + 1;
				
				write(mline, string'(" vo="));
				hwrite(mline, std_logic_vector(s_vo));
				writeline(output, mline);
			
			else
				s_enable <= '0';
			end if;
		
		end if;
		
	end process;

end behave;
